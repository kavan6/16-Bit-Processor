//Created by Kavan Heppenstall, 23/08/2003

module idecoder16bit(A, clk, );

endmodule