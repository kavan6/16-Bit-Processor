// Created by Kavan Heppenstall, 28/08/2024

module datapath();



endmodule